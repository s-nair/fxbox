library IEEE;
use IEEE.std_logic_1164.all;

-- Package Declaration Section
package fxbox_pkg is

	-- FXBOX TOP --

	constant MODE_COUNT_FX : natural := 3;
	constant CLK_TREE_LEN : natural := 15;
	
	
	-- DISPLAY DRIVER --
	
	constant CTR_LEN_DRV : natural := 10;
   
end package fxbox_pkg;

package body fxbox_pkg is
end package body fxbox_pkg;	